module python();

wire a;



endmodule