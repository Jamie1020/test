module python();
endmodule