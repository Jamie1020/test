module python();

wire a;
wire b;


endmodule